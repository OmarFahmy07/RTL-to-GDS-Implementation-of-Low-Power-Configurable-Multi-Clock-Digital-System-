module SYS_TOP_dft(input wire REF_CLK,
               input wire UART_CLK,
               input wire RST,
               input wire RX_IN,
               output wire TX_OUT,
               output wire PARITY_ERROR,
               output wire STOP_ERROR,
		// DFT Signals
	       input wire SI,
	       input wire SE,
	       input wire test_mode,
	       input wire scan_clk,
 	       input wire scan_rst,
	       output wire SO);
    
    //DFT Signals
    wire muxed_rst, muxed_rst1, muxed_rst2, muxed_ref_clk, muxed_uart_clk, muxed_uart_tx_clk;

    wire rst_sync_1_out;
    wire [7:0] RX_P_DATA;
    wire RX_D_VALID;
    wire RdData_Valid;
    wire Busy;
    wire [7:0] RdData;
    wire OUT_Valid;
    wire [15:0] ALU_OUT;
    wire [3:0] Address;
    wire [7:0] WrData;
    wire WrEn;
    wire RdEn;
    wire [3:0] ALU_FUN;
    wire ALU_EN;
    wire [7:0] TX_P_DATA;
    wire TX_D_VALID;
    wire CLK_EN;
    wire clk_div_en;
    wire [7:0] operand_A;
    wire [7:0] operand_B;
    wire [7:0] UART_config;
    wire [7:0] Div_ratio;
    wire ALU_CLK;
    wire TX_CLK;
    wire rst_sync_2_out;
    wire [7:0] P_DATA_TX;
    wire DATA_VALID_TX;
    wire BUSY_TX;
    wire [7:0] P_DATA_RX;
    wire DATA_VALID_RX;

    // Muxing ref clock
    mux2X1 U0_mux2X1 (
    .IN_0(REF_CLK),
    .IN_1(scan_clk),
    .sel(test_mode),
    .out(muxed_ref_clk)
    );

    // Muxing UART Rx clock
    mux2X1 U1_mux2X1 (
    .IN_0(UART_CLK),
    .IN_1(scan_clk),
    .sel(test_mode),
    .out(muxed_uart_clk)
    );

    // Muxing UART Tx clock
    mux2X1 U2_mux2X1 (
    .IN_0(TX_CLK),
    .IN_1(scan_clk),
    .sel(test_mode),
    .out(muxed_uart_tx_clk)
    );

    // Muxing reset 1
    mux2X1 U3_mux2X1 (
    .IN_0(rst_sync_1_out),
    .IN_1(scan_rst),
    .sel(test_mode),
    .out(muxed_rst1)
    );

    // Muxing reset 2
    mux2X1 U4_mux2X1 (
    .IN_0(rst_sync_2_out),
    .IN_1(scan_rst),
    .sel(test_mode),
    .out(muxed_rst2)
    );

    // Muxing reset
    mux2X1 U5_mux2X1 (
    .IN_0(RST),
    .IN_1(scan_rst),
    .sel(test_mode),
    .out(muxed_rst)
    );
    
    SYS_CTRL U0_SYS_CTRL
    (
    .clk(muxed_ref_clk),
    .rst(muxed_rst1),
    .RX_P_DATA(RX_P_DATA), // Rx data output
    .RX_D_VALID(RX_D_VALID), // Rx valid output
    .RdData_Valid(RdData_Valid), // Register file valid output
    .Busy(Busy), // Tx busy output
    .RdData(RdData), // Register file data output
    .OUT_Valid(OUT_Valid), // ALU valid output
    .ALU_OUT(ALU_OUT), // ALU data output
    .Address(Address), // Register file input address
    .WrData(WrData), // Register file input data
    .WrEn(WrEn), // Register file write enable
    .RdEn(RdEn), // Register file read enable
    .ALU_FUN(ALU_FUN), // ALU function selection
    .ALU_EN(ALU_EN), // ALU enable input
    .TX_P_DATA(TX_P_DATA), // Tx input data
    .TX_D_VALID(TX_D_VALID), // Tx input valid
    .CLK_EN(CLK_EN), // Clock gate enable
    .clk_div_en(clk_div_en) // Clock divider enable
    );
    
    Reg_File  #(.ADDRESS_WIDTH(4), .DATA_WIDTH(8)) U0_Reg_File
    (.WrEn(WrEn),
    .RdEn(RdEn),
    .Address(Address),
    .WrData(WrData),
    .CLK(muxed_ref_clk),
    .RST(muxed_rst1),
    .RdData(RdData),
    .RdData_Valid(RdData_Valid),
    .REG0(operand_A),
    .REG1(operand_B),
    .REG2(UART_config),
    .REG3(Div_ratio)
    );
    
    ALU #(.IN_DATA_WIDTH(8), .OUT_DATA_WIDTH(16)) U0_ALU
    (.A(operand_A),
    .B(operand_B),
    .func(ALU_FUN),
    .enable(ALU_EN),
    .clk(ALU_CLK),
    .rst(muxed_rst1),
    .result(ALU_OUT),
    .valid(OUT_Valid)
    );
    
    UART U0_UART
    (
    .TX_CLK(muxed_uart_tx_clk),
    .RX_CLK(muxed_uart_clk),
    .RST(muxed_rst2),
    .PAR_TYP(UART_config[1]),
    .PAR_EN(UART_config[0]),
    .P_DATA_TX(P_DATA_TX),
    .DATA_VALID_TX(DATA_VALID_TX),
    .RX_IN(RX_IN),
    .PRESCALE_RX(UART_config[7:2]),
    .TX_OUT(TX_OUT),
    .BUSY_TX(BUSY_TX),
    .P_DATA_RX(P_DATA_RX),
    .PAR_ERR_RX(PARITY_ERROR),
    .STP_ERR_RX(STOP_ERROR),
    .DATA_VALID_RX(DATA_VALID_RX)
    );
    
    CLK_GATE U0_CLK_GATE (
    .CLK_EN(CLK_EN | test_mode),
    .CLK(muxed_ref_clk),
    .GATED_CLK(ALU_CLK)
    );
    
    bit_synchronizer #(.BUS_WIDTH(1), .NUM_STAGES(2)) U0_bit_synchronizer
    (
    .ASYNC(BUSY_TX),
    .CLK(muxed_ref_clk),
    .RST(muxed_rst1),
    .SYNC(Busy)
    );
    
    data_synchronizer #(.BUS_WIDTH(8), .NUM_STAGES(2)) U0_data_sync_1
    (
    .unsync_bus(P_DATA_RX),
    .bus_enable(DATA_VALID_RX),
    .CLK(muxed_ref_clk),
    .RST(muxed_rst1),
    .sync_bus(RX_P_DATA),
    .enable_pulse(RX_D_VALID)
    );
    
    data_synchronizer #(.BUS_WIDTH(8), .NUM_STAGES(2)) U0_data_sync_2
    (
    .unsync_bus(TX_P_DATA),
    .bus_enable(TX_D_VALID),
    .CLK(muxed_uart_tx_clk),
    .RST(muxed_rst2),
    .sync_bus(P_DATA_TX),
    .enable_pulse(DATA_VALID_TX)
    );
    
    RST_SYNC #(.NUM_STAGES(2)) U0_RST_SYNC_1
    (
    .RST(muxed_rst),
    .CLK(muxed_ref_clk),
    .SYNC_RST(rst_sync_1_out)
    );
    
    RST_SYNC #(.NUM_STAGES(2)) U0_RST_SYNC_2
    (
    .RST(muxed_rst),
    .CLK(muxed_uart_clk),
    .SYNC_RST(rst_sync_2_out)
    );
    
    ClkDiv #(.RATIO_WIDTH(6)) U0_ClkDiv
    (.i_ref_clk(muxed_uart_clk),
    .i_rst_n(muxed_rst2),
    .i_clk_en(clk_div_en),
    .i_div_ratio(Div_ratio[5:0]),
    .o_div_clk(TX_CLK)
    );
    
endmodule
